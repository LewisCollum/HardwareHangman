library ieee, uart;
use ieee.std_logic_1164.all;

entity UARTAdapter is
  port(
    clock: in std_logic;
    reset: in std_logic);
end entity;

architecture behavioral of UARTAdapter is
begin

end architecture;
