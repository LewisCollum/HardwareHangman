package state_pkg is
  type PS2 is (ready, parse);
end package;
